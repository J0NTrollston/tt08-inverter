** sch_path: /home/ttuser/Documents/tt08-inverter/xschem/testbench.sch
**.subckt testbench in out
*.ipin in
*.opin out
x1 VSS net1 net2 in myInverter
V1 VSS GND 0
V2 VDD GND 1.8
R1 out net2 500 m=1
C1 net2 GND 5p m=1
Vmeas VDD net1 0
.save i(vmeas)
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.options savecurrents
vin in 0 pulse 0 1.8 5n 1n 1n 50n 100n
.control
save all
tran 100p 200n
write testbench.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  myInverter.sym # of pins=4
** sym_path: /home/ttuser/Documents/tt08-inverter/xschem/myInverter.sym
** sch_path: /home/ttuser/Documents/tt08-inverter/xschem/myInverter.sch
.subckt myInverter VSS VDD out in
*.iopin VDD
*.iopin VSS
*.ipin in
*.opin out
XM2 out in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
