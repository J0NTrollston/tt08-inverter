magic
tech sky130A
magscale 1 2
timestamp 1726789828
<< pwell >>
rect 1096 -1852 1374 -1794
<< viali >>
rect 1272 286 1402 322
rect 1274 -1938 1400 -1904
<< metal1 >>
rect -122 784 1650 984
rect 725 126 923 784
rect 1261 322 1416 784
rect 1261 286 1272 322
rect 1402 286 1416 322
rect 1261 273 1416 286
rect 979 175 985 237
rect 1047 236 1107 237
rect 1047 178 1372 236
rect 1047 175 1107 178
rect 637 -249 1311 126
rect 1365 44 2089 125
rect 1365 -156 2384 44
rect 1365 -237 2089 -156
rect 979 -360 985 -298
rect 1047 -360 1374 -298
rect 980 -728 1042 -360
rect -122 -928 1042 -728
rect 980 -1473 1042 -928
rect 2184 -730 2384 -156
rect 2184 -930 3172 -730
rect 979 -1531 985 -1473
rect 1043 -1474 1103 -1473
rect 1043 -1531 1374 -1474
rect 1058 -1534 1374 -1531
rect 734 -1763 1312 -1562
rect 2190 -1566 2390 -930
rect 1870 -1580 2390 -1566
rect 1367 -1751 2390 -1580
rect 734 -2101 935 -1763
rect 1870 -1766 2390 -1751
rect 979 -1852 985 -1794
rect 1043 -1852 1374 -1794
rect 1239 -1904 1440 -1888
rect 1239 -1938 1274 -1904
rect 1400 -1938 1440 -1904
rect 1239 -2101 1440 -1938
rect -122 -2302 1656 -2101
<< via1 >>
rect 985 175 1047 237
rect 985 -360 1047 -298
rect 985 -1531 1043 -1473
rect 985 -1852 1043 -1794
<< metal2 >>
rect 985 237 1047 243
rect 985 -298 1047 175
rect 985 -366 1047 -360
rect 985 -1473 1043 -1467
rect 985 -1794 1043 -1531
rect 985 -1858 1043 -1852
use sky130_fd_pr__pfet_01v8_XGAKDL  XM1
timestamp 1726789828
transform 1 0 1339 0 1 -61
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1726789828
transform 1 0 1339 0 1 -1664
box -211 -310 211 310
<< labels >>
flabel metal1 -122 -928 78 -728 0 FreeSans 256 0 0 0 in
port 3 nsew
flabel metal1 -122 -2302 78 -2102 0 FreeSans 256 0 0 0 VSS
port 0 nsew
flabel metal1 -122 784 78 984 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 2972 -930 3172 -730 0 FreeSans 256 0 0 0 out
port 2 nsew
<< end >>
