** sch_path: /home/ttuser/Documents/tt08-inverter/xschem/myInverter.sch
.subckt myInverter VSS VDD out in
*.PININFO VDD:B VSS:B in:I out:O
XM2 out in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM1 out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
.ends
.end
